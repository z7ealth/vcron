module types

pub struct Cron {
	minutes u8
	hours u8
	days u8
	month u8
	week_days u8
}